package parameters;

// Specific configuration bus size parameters
typedef 8 CBADDRSIZE;  //size of configuration address bus to decode
typedef 16 CBDATASIZE; //size of configuration data bus 

endpackage
