package parameters;

typedef 8 CBADDRSIZE;  //size of configuration address bus to decode
// Change the below line to generate the K-bit integer Matrix adder (currently it is 16-bit integer Matrix adder)
typedef 16 CBDATASIZE; //size of configuration data bus and the register used in the Accelerator

endpackage
